magic
tech sky130A
magscale 1 2
timestamp 1769561617
<< nwell >>
rect -308 -418 308 418
<< mvpmos >>
rect -50 -121 50 121
<< mvpdiff >>
rect -108 109 -50 121
rect -108 -109 -96 109
rect -62 -109 -50 109
rect -108 -121 -50 -109
rect 50 109 108 121
rect 50 -109 62 109
rect 96 -109 108 109
rect 50 -121 108 -109
<< mvpdiffc >>
rect -96 -109 -62 109
rect 62 -109 96 109
<< mvnsubdiff >>
rect -242 340 242 352
rect -242 306 -134 340
rect 134 306 242 340
rect -242 294 242 306
rect -242 244 -184 294
rect -242 -244 -230 244
rect -196 -244 -184 244
rect 184 244 242 294
rect -242 -294 -184 -244
rect 184 -244 196 244
rect 230 -244 242 244
rect 184 -294 242 -244
rect -242 -306 242 -294
rect -242 -340 -134 -306
rect 134 -340 242 -306
rect -242 -352 242 -340
<< mvnsubdiffcont >>
rect -134 306 134 340
rect -230 -244 -196 244
rect 196 -244 230 244
rect -134 -340 134 -306
<< poly >>
rect -50 202 50 218
rect -50 168 -34 202
rect 34 168 50 202
rect -50 121 50 168
rect -50 -168 50 -121
rect -50 -202 -34 -168
rect 34 -202 50 -168
rect -50 -218 50 -202
<< polycont >>
rect -34 168 34 202
rect -34 -202 34 -168
<< locali >>
rect -230 306 -134 340
rect 134 306 230 340
rect -230 244 -196 306
rect 196 244 230 306
rect -50 168 -34 202
rect 34 168 50 202
rect -96 109 -62 125
rect -96 -125 -62 -109
rect 62 109 96 125
rect 62 -125 96 -109
rect -50 -202 -34 -168
rect 34 -202 50 -168
rect -230 -306 -196 -244
rect 196 -306 230 -244
rect -230 -340 -134 -306
rect 134 -340 230 -306
<< viali >>
rect -34 168 34 202
rect -96 -109 -62 109
rect 62 -109 96 109
rect -34 -202 34 -168
<< metal1 >>
rect -46 202 46 208
rect -46 168 -34 202
rect 34 168 46 202
rect -46 162 46 168
rect -102 109 -56 121
rect -102 -109 -96 109
rect -62 -109 -56 109
rect -102 -121 -56 -109
rect 56 109 102 121
rect 56 -109 62 109
rect 96 -109 102 109
rect 56 -121 102 -109
rect -46 -168 46 -162
rect -46 -202 -34 -168
rect 34 -202 46 -168
rect -46 -208 46 -202
<< properties >>
string FIXED_BBOX -213 -323 213 323
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1.21 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
