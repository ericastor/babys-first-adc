magic
tech sky130A
magscale 1 2
timestamp 1769561617
<< pwell >>
rect -278 -383 278 383
<< mvnmos >>
rect -50 -125 50 125
<< mvndiff >>
rect -108 113 -50 125
rect -108 -113 -96 113
rect -62 -113 -50 113
rect -108 -125 -50 -113
rect 50 113 108 125
rect 50 -113 62 113
rect 96 -113 108 113
rect 50 -125 108 -113
<< mvndiffc >>
rect -96 -113 -62 113
rect 62 -113 96 113
<< mvpsubdiff >>
rect -242 335 242 347
rect -242 301 -134 335
rect 134 301 242 335
rect -242 289 242 301
rect -242 239 -184 289
rect -242 -239 -230 239
rect -196 -239 -184 239
rect 184 239 242 289
rect -242 -289 -184 -239
rect 184 -239 196 239
rect 230 -239 242 239
rect 184 -289 242 -239
rect -242 -301 242 -289
rect -242 -335 -134 -301
rect 134 -335 242 -301
rect -242 -347 242 -335
<< mvpsubdiffcont >>
rect -134 301 134 335
rect -230 -239 -196 239
rect 196 -239 230 239
rect -134 -335 134 -301
<< poly >>
rect -50 197 50 213
rect -50 163 -34 197
rect 34 163 50 197
rect -50 125 50 163
rect -50 -163 50 -125
rect -50 -197 -34 -163
rect 34 -197 50 -163
rect -50 -213 50 -197
<< polycont >>
rect -34 163 34 197
rect -34 -197 34 -163
<< locali >>
rect -230 301 -134 335
rect 134 301 230 335
rect -230 239 -196 301
rect 196 239 230 301
rect -50 163 -34 197
rect 34 163 50 197
rect -96 113 -62 129
rect -96 -129 -62 -113
rect 62 113 96 129
rect 62 -129 96 -113
rect -50 -197 -34 -163
rect 34 -197 50 -163
rect -230 -301 -196 -239
rect 196 -301 230 -239
rect -230 -335 -134 -301
rect 134 -335 230 -301
<< viali >>
rect -34 163 34 197
rect -96 -113 -62 113
rect 62 -113 96 113
rect -34 -197 34 -163
<< metal1 >>
rect -46 197 46 203
rect -46 163 -34 197
rect 34 163 46 197
rect -46 157 46 163
rect -102 113 -56 125
rect -102 -113 -96 113
rect -62 -113 -56 113
rect -102 -125 -56 -113
rect 56 113 102 125
rect 56 -113 62 113
rect 96 -113 102 113
rect 56 -125 102 -113
rect -46 -163 46 -157
rect -46 -197 -34 -163
rect 34 -197 46 -163
rect -46 -203 46 -197
<< properties >>
string FIXED_BBOX -213 -318 213 318
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1.25 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
