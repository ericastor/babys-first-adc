magic
tech sky130A
magscale 1 2
timestamp 1769561617
<< metal3 >>
rect -1986 1812 1986 1840
rect -1986 -1812 1902 1812
rect 1966 -1812 1986 1812
rect -1986 -1840 1986 -1812
<< via3 >>
rect 1902 -1812 1966 1812
<< mimcap >>
rect -1946 1760 1654 1800
rect -1946 -1760 -1906 1760
rect 1614 -1760 1654 1760
rect -1946 -1800 1654 -1760
<< mimcapcontact >>
rect -1906 -1760 1614 1760
<< metal4 >>
rect 1886 1812 1982 1828
rect -1907 1760 1615 1761
rect -1907 -1760 -1906 1760
rect 1614 -1760 1615 1760
rect -1907 -1761 1615 -1760
rect 1886 -1812 1902 1812
rect 1966 -1812 1982 1812
rect 1886 -1828 1982 -1812
<< properties >>
string FIXED_BBOX -1986 -1840 1694 1840
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 18.0 l 18.0 val 661.68 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
