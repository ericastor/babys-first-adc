** sch_path: /home/ttuser/babys-first-adc/xschem/track_testbench.sch
**.subckt track_testbench out
*.opin out
VDD_src VDD GND 3.3
VSS_src VSS GND 0
V4 in VSS 0 ac 1 0 sin(1.65 1.65 33e6 0 0 0)
XM1 VDD out net1 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
R1 net1 VSS 1 m=1
Vclk CLK VSS 0
Vclk1 CLKB VSS 3.3
x1 CLK CLKB VDD VSS out in track_and_hold
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/ttuser/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt





  .option savecurrents
  .control
    tran 0.05n 3u
    remzerovec
    write track_testbench.raw

    let in_spec = in - 1.65
    let out_spec = out - 1.65
    linearize in_spec out_spec
    fft in_spec out_spec
    set appendwrite
    write track_testbench.raw
  .endc



**** end user architecture code
**.ends

* expanding   symbol:  track_and_hold.sym # of pins=6
** sym_path: /home/ttuser/babys-first-adc/xschem/track_and_hold.sym
** sch_path: /home/ttuser/babys-first-adc/xschem/track_and_hold.sch
.subckt track_and_hold HLD TRK VDD VSS out in
*.iopin VSS
*.iopin VDD
*.ipin in
*.opin out
*.iopin TRK
*.iopin HLD
XC1 out VSS sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=1 m=1
V1 net2 in 3.3
XM1 out net1 in VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
R1 VDD VSS 1G m=1
S2 net1 net2 TRK VSS SWITCH1
S4 net1 VSS HLD VSS SWITCH1
**** begin user architecture code



.model switch1 sw vt=1.65 vh=0 ron=1 roff=1G



**** end user architecture code
V2 in net3 3.3
S2p net4 net3 TRK VSS SWITCH1
S4p net4 VDD HLD VSS SWITCH1
XM2 out net4 in VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1.36 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
