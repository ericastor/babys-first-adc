** sch_path: /home/ttuser/babys-first-adc/xschem/testbench.sch
**.subckt testbench out
*.opin out
VDD_src VDD GND 3.3
VSS_src VSS GND 0
V4 in VSS 0 ac 1 0 sin(1.65 1.65 7e6 0 0 90)
XM1 net2 out net1 GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
R1 net1 GND 1 m=1
Vclk CLK VSS 0 ac 1 0 pulse(3.3 0 0 0.1ns 0.1ns 7.5ns 15ns)
Vclk1 CLKB VSS 0 ac 1 0 pulse(0 3.3 0 0.1ns 0.1ns 7.5ns 15ns)
x1 CLK CLKB VDD VSS out in parametric_track_and_hold WT=1 PFT=1.21 PF=2 WS=5 WB=5 CB=18
V_test net2 GND 3.3
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/ttuser/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt





  .option savecurrents
  .control
    tran 0.05n 6u
    remzerovec
    write testbench.raw

    let lin-tstart = 12.5n
    let lin-tstep = 15n
    let in_spec = in - 1.65
    let out_spec = out - 1.65
    linearize in_spec out_spec
    fft in_spec out_spec
    set appendwrite
    write testbench.raw

    meas sp peak_noise MAX vdb(out_spec) from=1Meg to=6Meg
    echo "Peak noise < 6Meg: $&peak_noise dB"

    meas sp peak_harmonic MAX vdb(out_spec) from=10Meg to=33Meg
    echo "Peak harmonic: $&peak_harmonic dB"

    setplot tran1
    let s = (VDD_src#branch)^2
    meas tran ms AVG s
    let rms = 1000*sqrt(ms)
    echo "RMS current (from VDD): $&rms mA"
  .endc



**** end user architecture code
**.ends

* expanding   symbol:  parametric_track_and_hold.sym # of pins=6
** sym_path: /home/ttuser/babys-first-adc/xschem/parametric_track_and_hold.sym
** sch_path: /home/ttuser/babys-first-adc/xschem/parametric_track_and_hold.sch
.subckt parametric_track_and_hold HLD TRK VDD VSS out in  WT=1 PFT=1.21 PF=2 WS=5 WB=5 CB=18
*.iopin VSS
*.iopin VDD
*.ipin in
*.opin out
*.iopin HLD
*.iopin TRK
XC2 out VSS sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=1 m=1
XM1 out X in VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W={WT} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1p out Xp in VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W={WT*PFT} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 net1 HLD VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W={2*WS} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 P Y X P sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W={WS*PF} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 in X Q VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W={WB} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 Q HLD VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W={WB} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3p Qp Xp in VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W={WB*PF} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 P X VDD P sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W={WB*PF} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XCb P Q sky130_fd_pr__cap_mim_m3_1 W={CB} L={CB} MF=1 m=1
XM8 X VDD net1 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W={2*WS} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMb Y TRK VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W={(WS/4)*PF} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMa Y TRK Q VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W={WS/10} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMc Q X Y VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W={WS} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XCbp Pp Qp sky130_fd_pr__cap_mim_m3_1 W={CB} L={CB} MF=1 m=1
XM6p VDD TRK Qp VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W={WB*PF} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5p VSS Xp Pp Pp sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W={WB} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2p Xp net2 Pp Pp sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W={WS} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMcp net2 Xp Qp VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W={WS*PF} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMap Qp HLD net2 VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W={(WS/10)*PF} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMbp VSS HLD net2 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W={WS/4} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8p net3 VSS Xp VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W={2*WS*PF} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4p VDD TRK net3 VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W={2*WS*PF} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
