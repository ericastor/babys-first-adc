magic
tech sky130A
timestamp 1769561617
<< pwell >>
rect -139 -154 139 154
<< mvnmos >>
rect -25 -25 25 25
<< mvndiff >>
rect -54 19 -25 25
rect -54 -19 -48 19
rect -31 -19 -25 19
rect -54 -25 -25 -19
rect 25 19 54 25
rect 25 -19 31 19
rect 48 -19 54 19
rect 25 -25 54 -19
<< mvndiffc >>
rect -48 -19 -31 19
rect 31 -19 48 19
<< mvpsubdiff >>
rect -121 130 121 136
rect -121 113 -67 130
rect 67 113 121 130
rect -121 107 121 113
rect -121 82 -92 107
rect -121 -82 -115 82
rect -98 -82 -92 82
rect 92 82 121 107
rect -121 -107 -92 -82
rect 92 -82 98 82
rect 115 -82 121 82
rect 92 -107 121 -82
rect -121 -113 121 -107
rect -121 -130 -67 -113
rect 67 -130 121 -113
rect -121 -136 121 -130
<< mvpsubdiffcont >>
rect -67 113 67 130
rect -115 -82 -98 82
rect 98 -82 115 82
rect -67 -130 67 -113
<< poly >>
rect -25 61 25 69
rect -25 44 -17 61
rect 17 44 25 61
rect -25 25 25 44
rect -25 -44 25 -25
rect -25 -61 -17 -44
rect 17 -61 25 -44
rect -25 -69 25 -61
<< polycont >>
rect -17 44 17 61
rect -17 -61 17 -44
<< locali >>
rect -115 113 -67 130
rect 67 113 115 130
rect -115 82 -98 113
rect 98 82 115 113
rect -25 44 -17 61
rect 17 44 25 61
rect -48 19 -31 27
rect -48 -27 -31 -19
rect 31 19 48 27
rect 31 -27 48 -19
rect -25 -61 -17 -44
rect 17 -61 25 -44
rect -115 -113 -98 -82
rect 98 -113 115 -82
rect -115 -130 -67 -113
rect 67 -130 115 -113
<< viali >>
rect -17 44 17 61
rect -48 -19 -31 19
rect 31 -19 48 19
rect -17 -61 17 -44
<< metal1 >>
rect -23 61 23 64
rect -23 44 -17 61
rect 17 44 23 61
rect -23 41 23 44
rect -51 19 -28 25
rect -51 -19 -48 19
rect -31 -19 -28 19
rect -51 -25 -28 -19
rect 28 19 51 25
rect 28 -19 31 19
rect 48 -19 51 19
rect 28 -25 51 -19
rect -23 -44 23 -41
rect -23 -61 -17 -44
rect 17 -61 23 -44
rect -23 -64 23 -61
<< properties >>
string FIXED_BBOX -106 -121 106 121
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 0.5 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
