** sch_path: /home/ttuser/babys-first-adc/xschem/track_and_hold.sch
.subckt track_and_hold HLD TRK VDD VSS out in
*.PININFO VSS:B VDD:B in:I out:O HLD:B TRK:B
XC1 out VSS sky130_fd_pr__cap_mim_m3_1 W=5 L=5 m=1
XM1 out X in VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM1p out Xp in VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1.21 nf=1 m=1
XM4 net1 HLD VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 nf=1 m=1
XM2 P Y X P sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=10 nf=1 m=1
XM3 in X Q VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 nf=1 m=1
XM6 Q HLD VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 nf=1 m=1
XM3p Qp Xp in VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=10 nf=1 m=1
XM5 P X VDD P sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=10 nf=1 m=1
XCb P Q sky130_fd_pr__cap_mim_m3_1 W=18 L=18 m=1
XM8 X VDD net1 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 nf=1 m=1
XMb Y TRK VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2.5 nf=1 m=1
XMa Y TRK Q VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.5 nf=1 m=1
XMc Q X Y VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 nf=1 m=1
XCbp Pp Qp sky130_fd_pr__cap_mim_m3_1 W=18 L=18 m=1
XM6p VDD TRK Qp VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=10 nf=1 m=1
XM5p VSS Xp Pp Pp sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 nf=1 m=1
XM2p Xp Yp Pp Pp sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 nf=1 m=1
XMcp Yp Xp Qp VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=10 nf=1 m=1
XMap Qp HLD Yp VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XMbp VSS HLD Yp VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.25 nf=1 m=1
XM8p net2 VSS Xp VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=20 nf=1 m=1
XM4p VDD TRK net2 VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=20 nf=1 m=1
.ends
.end
