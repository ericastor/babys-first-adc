** sch_path: /home/ttuser/babys-first-adc/xschem/sample_and_hold.sch
**.subckt sample_and_hold VDD VSS HLD TRK out in
*.iopin VSS
*.iopin VDD
*.ipin in
*.opin out
*.iopin TRK
*.iopin HLD
XC1 out VSS sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
V1 net1 in 3.3
XM1 out gate in VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
R1 VDD VSS 1G m=1
S1 gate net1 TRK VSS SWITCH1
S2 gate VSS HLD VSS SWITCH1
V2 in net2 3.3
S3 net3 net2 TRK VSS SWITCH1
S4 net3 VDD HLD VSS SWITCH1
XM2 out net3 in VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code



.model switch1 sw vt=1.65 vh=0 ron=1 roff=1G



**** end user architecture code
**.ends
.end
