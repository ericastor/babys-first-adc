** sch_path: /home/ttuser/babys-first-adc/xschem/hold_testbench.sch
**.subckt hold_testbench out
*.opin out
VDD_src VDD GND 3.3
VSS_src VSS GND 0
V4 in VSS 3
XM1 VDD out net1 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
R1 net1 VSS 1 m=1
Vclk TRK VSS 0 ac 1 0 pulse(3.3 0 0 0.1ns 0.1ns 50ns 100ns)
Vclk1 HLD VSS 0 ac 1 0 pulse(0 3.3 0 0.1ns 0.1ns 50ns 100ns)
x1 HLD TRK VDD VSS out in parametric_track_and_hold WT=1 PFT=1.21 PF=2 WS=5 WB=5 CB=18
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/ttuser/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice ss





.control
  let v_start = 0
  let v_stop  = 3.3
  let v_step  = 0.1
  let n_points = floor((v_stop - v_start) / v_step) + 1

  let index = 0

  * Initialize vectors in the 'const' plot
  let in_vec = v_start + (v_stop - v_start) * vector(n_points) / (n_points - 1)
  let diff_vec = vector($&n_points)

  set temp=27

  while $&index < $&n_points
    destroy all

    alter V4 = in_vec[$&index]
    tran 0.1n 110n

    meas tran v_prehold find v(out) at=95n
    meas tran v_earlyhold find v(out) at=105n

    let d_val = v_earlyhold - v_prehold
    let const.diff_vec[index] = d_val

    let index = index + 1
  end

  let v_tracked = const.in_vec
  let hold_delta = const.diff_vec

  setscale v_tracked hold_delta
  settype voltage v_tracked hold_delta
  plot hold_delta vs v_tracked
  let v = v_tracked[0]
  let d = hold_delta[0] * 1000
  echo "$&d mV \@ $&v V"
  let v = v_tracked[$&n_points - 1]
  let d = hold_delta[$&n_points - 1] * 1000
  echo "$&d mV \@ $&v V"
.endc



**** end user architecture code
**.ends

* expanding   symbol:  parametric_track_and_hold.sym # of pins=6
** sym_path: /home/ttuser/babys-first-adc/xschem/parametric_track_and_hold.sym
** sch_path: /home/ttuser/babys-first-adc/xschem/parametric_track_and_hold.sch
.subckt parametric_track_and_hold HLD TRK VDD VSS out in  WT=1 PFT=1.21 PF=2 WS=5 WB=5 CB=18
*.iopin VSS
*.iopin VDD
*.ipin in
*.opin out
*.iopin TRK
*.iopin HLD
XC1 out VSS sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=1 m=1
XM1 out X in VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W={WT} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1p out net1 in VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W={WT*PFT} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 VSS HLD X VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W={WS} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4p net1 TRK VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W={WS*PF} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 X HLD P P sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W={WS*PF} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2p net2 TRK net1 net2 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W={WS} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 in X Q VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W={WB} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 Q HLD VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W={WB} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3p net3 net1 in VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W={WB*PF} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6p VDD TRK net3 VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W={WB*PF} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 P X VDD P sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W={WB*PF} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XCb P Q sky130_fd_pr__cap_mim_m3_1 W={CB} L={CB} MF=1 m=1
XCbp net2 net3 sky130_fd_pr__cap_mim_m3_1 W={CB} L={CB} MF=1 m=1
XM5p VSS net1 net2 net2 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W={WB*PF} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
