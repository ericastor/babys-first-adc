magic
tech sky130A
magscale 1 2
timestamp 1769749962
<< dnwell >>
rect 5820 -2340 7520 -220
<< nwell >>
rect 1300 -1000 1740 -400
rect 5920 -520 7420 -320
rect 1300 -1620 1560 -1000
rect 5920 -2040 6120 -520
rect 7220 -2040 7420 -520
rect 5920 -2240 7420 -2040
rect 840 -3020 1480 -2980
<< nsubdiff >>
rect 5960 -380 7380 -360
rect 5960 -400 6020 -380
rect 7340 -400 7380 -380
rect 5960 -2160 5980 -400
rect 6060 -480 7280 -460
rect 6060 -2080 6080 -480
rect 7260 -2080 7280 -480
rect 6060 -2100 7280 -2080
rect 7360 -2160 7380 -400
rect 5960 -2180 6000 -2160
rect 7340 -2180 7380 -2160
rect 5960 -2200 7380 -2180
<< nsubdiffcont >>
rect 6020 -400 7340 -380
rect 5980 -460 7360 -400
rect 5980 -2100 6060 -460
rect 7280 -2100 7360 -460
rect 5980 -2160 7360 -2100
rect 6000 -2180 7340 -2160
<< locali >>
rect 5960 -380 7380 -360
rect 5960 -400 6020 -380
rect 7340 -400 7380 -380
rect 5960 -2160 5980 -400
rect 6060 -480 7280 -460
rect 6060 -2080 6080 -480
rect 7260 -2080 7280 -480
rect 6060 -2100 7280 -2080
rect 7360 -2160 7380 -400
rect 5960 -2180 6000 -2160
rect 7340 -2180 7380 -2160
rect 5960 -2200 7380 -2180
<< viali >>
rect 3320 3640 3360 3680
rect 3320 3540 3360 3580
rect 3600 2460 3640 2520
rect 3600 2280 3640 2340
rect 3260 920 3300 960
rect 3400 920 3440 960
rect 1640 880 1680 920
rect 3320 800 3360 840
rect 4780 620 4820 660
rect 1040 500 1080 540
rect 940 -520 980 -480
rect 1780 -520 1820 -480
rect 4380 -920 4420 -880
rect 2200 -1320 2240 -1280
rect 2380 -1320 2420 -1280
rect 5980 -1080 6060 -920
rect 6580 -1300 6640 -1260
rect 6700 -1300 6760 -1260
rect 1900 -2330 1940 -2290
rect 3020 -3120 3060 -3080
rect 3020 -4140 3060 -4100
<< metal1 >>
rect 3234 4140 3240 4160
rect 2620 3960 3240 4140
rect 3440 4140 3446 4160
rect 3440 3960 4600 4140
rect 2620 3940 4600 3960
rect 2280 3920 2360 3926
rect 0 3700 560 3900
rect 2360 3900 2580 3920
rect 2360 3860 4660 3900
rect 2360 3840 2580 3860
rect 2280 3834 2360 3840
rect 2620 3740 4600 3820
rect 360 3440 560 3700
rect 3300 3680 3380 3700
rect 3300 3640 3320 3680
rect 3360 3640 3380 3680
rect 3294 3560 3300 3640
rect 3380 3560 3386 3640
rect 3300 3540 3320 3560
rect 3360 3540 3380 3560
rect 3300 3520 3380 3540
rect 4520 3480 4600 3740
rect 360 3240 1580 3440
rect 1780 3360 2560 3440
rect 2620 3400 4600 3480
rect 1780 3320 4660 3360
rect 1780 3240 2560 3320
rect 2240 3160 2440 3240
rect 2620 3200 4600 3280
rect 2240 2960 2800 3160
rect 4520 3100 4600 3200
rect 4520 3020 4840 3100
rect 2600 2760 4600 2960
rect 4760 2740 4840 3020
rect 4640 2720 4840 2740
rect 2540 2680 4840 2720
rect 4640 2660 4840 2680
rect 2600 2560 4580 2640
rect 3580 2520 3660 2560
rect 3580 2460 3600 2520
rect 3640 2460 3660 2520
rect 3580 2440 3660 2460
rect 3580 2340 3660 2360
rect 3580 2280 3600 2340
rect 3640 2280 3660 2340
rect 3580 2240 3660 2280
rect 2620 2160 4580 2240
rect 2480 2120 2560 2140
rect 0 2040 200 2100
rect 2480 2080 4660 2120
rect 1160 2040 1240 2046
rect 0 1960 1160 2040
rect 0 1900 200 1960
rect 1160 1740 1240 1960
rect 1060 780 1140 1700
rect 1020 700 1140 780
rect 1020 540 1100 700
rect 1180 640 1220 1740
rect 1260 780 1340 1700
rect 2480 1320 2560 2080
rect 2600 1960 4600 2040
rect 4520 1800 4600 1960
rect 4760 1800 4840 2660
rect 4520 1720 4840 1800
rect 2260 1280 3700 1320
rect 2260 1240 4600 1280
rect 1860 1160 2340 1240
rect 3620 1200 4600 1240
rect 2660 1160 2960 1180
rect 4640 1160 4720 1720
rect 2420 1120 2660 1140
rect 1780 1080 2660 1120
rect 2740 1120 3160 1160
rect 3540 1120 4720 1160
rect 2740 1100 2960 1120
rect 2420 1060 2740 1080
rect 1840 980 2360 1040
rect 1580 940 2360 980
rect 1580 860 1620 940
rect 1740 860 2360 940
rect 1580 820 2360 860
rect 3000 780 3100 1080
rect 3600 1000 4600 1080
rect 3240 960 3300 980
rect 3240 920 3260 960
rect 3240 900 3300 920
rect 3380 960 3460 980
rect 3380 920 3400 960
rect 3440 920 3460 960
rect 3380 900 3460 920
rect 3300 840 3380 900
rect 3300 800 3320 840
rect 3360 800 3380 840
rect 3300 780 3380 800
rect 1340 740 3100 780
rect 3920 740 4000 1000
rect 1340 700 4000 740
rect 1260 694 1340 700
rect 3000 660 4000 700
rect 4640 640 4720 1120
rect 7400 940 7600 1000
rect 5560 860 7600 940
rect 4060 620 4720 640
rect 2940 580 4720 620
rect 4754 600 4760 680
rect 4840 600 4846 680
rect 4060 560 4720 580
rect 1020 500 1040 540
rect 1080 500 1100 540
rect 3940 500 4000 540
rect 4540 500 4660 560
rect 1020 306 1100 500
rect 3000 460 4000 500
rect 3920 400 4540 460
rect 980 300 1180 306
rect 1180 100 2800 300
rect 3000 100 3006 300
rect 4420 260 4540 400
rect 0 40 200 100
rect 980 94 1180 100
rect 4420 40 4500 260
rect 4580 200 4620 500
rect 4700 340 4740 460
rect 4700 300 4780 340
rect 4660 260 4780 300
rect 0 -40 4500 40
rect 0 -100 200 -40
rect 920 -460 1840 -400
rect 920 -480 1760 -460
rect 920 -520 940 -480
rect 980 -520 1760 -480
rect 4420 -460 4500 -40
rect 4700 40 4780 260
rect 5560 60 5640 860
rect 7400 800 7600 860
rect 5540 40 5660 60
rect 4700 -40 5560 40
rect 5640 -40 5660 40
rect 4420 -520 4540 -460
rect 920 -700 1040 -520
rect 1760 -546 1840 -540
rect 3920 -560 4540 -520
rect 2000 -600 4540 -560
rect 3940 -640 4000 -600
rect 920 -760 1100 -700
rect 960 -2700 1100 -760
rect 0 -2740 200 -2700
rect 1140 -2734 1180 -640
rect 4060 -680 4340 -660
rect 1940 -720 4340 -680
rect 4500 -700 4540 -600
rect 4060 -740 4340 -720
rect 4580 -740 4620 -400
rect 4700 -460 4780 -40
rect 5540 -60 5660 -40
rect 4660 -500 4780 -460
rect 4700 -560 4780 -500
rect 4700 -700 4740 -560
rect 6220 -620 6980 -540
rect 1220 -960 1300 -954
rect 2000 -960 2040 -760
rect 1300 -1040 2040 -960
rect 1220 -1046 1300 -1040
rect 2000 -1160 2040 -1040
rect 2214 -1100 2220 -900
rect 2420 -1100 2960 -900
rect 3160 -1100 3166 -900
rect 1980 -1180 2040 -1160
rect 1960 -1200 2040 -1180
rect 1960 -1240 2020 -1200
rect 3960 -1240 4000 -760
rect 4260 -820 4720 -740
rect 4354 -940 4360 -860
rect 4440 -940 4446 -860
rect 1700 -1280 1760 -1260
rect 2180 -1280 2280 -1260
rect 1700 -1320 2080 -1280
rect 2180 -1320 2200 -1280
rect 2240 -1320 2280 -1280
rect 1700 -1680 1760 -1320
rect 2180 -1340 2280 -1320
rect 2360 -1280 2440 -1260
rect 4640 -1280 4720 -820
rect 6220 -780 6300 -620
rect 6220 -860 6340 -780
rect 5920 -900 6120 -894
rect 5920 -1106 6120 -1100
rect 2360 -1320 2380 -1280
rect 2420 -1320 2440 -1280
rect 2540 -1320 4720 -1280
rect 2360 -1340 2440 -1320
rect 1820 -1440 2020 -1360
rect 2600 -1440 4600 -1360
rect 1574 -1760 1580 -1680
rect 1660 -1760 1760 -1680
rect 1680 -2080 1760 -1760
rect 1880 -1740 1960 -1440
rect 3480 -1740 3560 -1440
rect 4640 -1620 4720 -1320
rect 6260 -1620 6340 -860
rect 4640 -1700 6340 -1620
rect 1880 -1820 3560 -1740
rect 1880 -1960 1960 -1820
rect 3480 -1940 3560 -1820
rect 1800 -2040 2040 -1960
rect 3480 -2026 3560 -2020
rect 1680 -2120 2100 -2080
rect 1680 -2140 1760 -2120
rect 1800 -2240 2040 -2160
rect 1820 -2290 2020 -2240
rect 1820 -2320 1900 -2290
rect 1940 -2320 2020 -2290
rect 2020 -2520 3380 -2320
rect 1820 -2526 2020 -2520
rect 1120 -2740 1200 -2734
rect 0 -2820 1120 -2740
rect 0 -2900 200 -2820
rect 1120 -2826 1200 -2820
rect 3180 -2740 3380 -2520
rect 4400 -2740 4600 -2734
rect 3180 -2940 4400 -2740
rect 4400 -2946 4600 -2940
rect 2994 -3140 3000 -3060
rect 3080 -3140 3086 -3060
rect 4740 -3180 4820 -1700
rect 6260 -1780 6340 -1700
rect 6380 -1820 6420 -720
rect 6900 -740 6980 -620
rect 6460 -1260 6880 -780
rect 6460 -1300 6580 -1260
rect 6640 -1300 6700 -1260
rect 6760 -1300 6880 -1260
rect 6460 -1660 6880 -1300
rect 6460 -1760 6620 -1660
rect 6720 -1760 6880 -1660
rect 6460 -1780 6880 -1760
rect 6354 -1900 6360 -1820
rect 6440 -1900 6446 -1820
rect 6920 -1840 6960 -740
rect 7000 -1680 7080 -780
rect 7000 -1780 7120 -1680
rect 7040 -2740 7120 -1780
rect 4960 -2760 7120 -2740
rect 4960 -2920 4980 -2760
rect 5140 -2920 7120 -2760
rect 4960 -2940 7120 -2920
rect 360 -3220 560 -3214
rect 560 -3290 850 -3230
rect 900 -3260 4900 -3180
rect 560 -3330 4950 -3290
rect 560 -3390 850 -3330
rect 360 -3700 560 -3420
rect 920 -3440 4880 -3380
rect 0 -3900 560 -3700
rect 4740 -3780 4820 -3440
rect 920 -3840 4880 -3780
rect 760 -3870 860 -3860
rect 760 -3950 780 -3870
rect 860 -3890 866 -3870
rect 860 -3930 4950 -3890
rect 860 -3950 866 -3930
rect 760 -3960 860 -3950
rect 2960 -3980 3000 -3960
rect 920 -4180 3000 -3980
rect 3120 -3980 3160 -3960
rect 3120 -4180 4880 -3980
rect 920 -4220 4880 -4180
<< via1 >>
rect 3240 3960 3440 4160
rect 2280 3840 2360 3920
rect 3300 3580 3380 3640
rect 3300 3560 3320 3580
rect 3320 3560 3360 3580
rect 3360 3560 3380 3580
rect 1580 3240 1780 3440
rect 3580 2360 3660 2440
rect 1160 1960 1240 2040
rect 2660 1080 2740 1160
rect 1620 920 1740 940
rect 1620 880 1640 920
rect 1640 880 1680 920
rect 1680 880 1740 920
rect 1620 860 1740 880
rect 3300 900 3380 980
rect 1260 700 1340 780
rect 4760 660 4840 680
rect 4760 620 4780 660
rect 4780 620 4820 660
rect 4820 620 4840 660
rect 4760 600 4840 620
rect 980 100 1180 300
rect 2800 100 3000 300
rect 1760 -480 1840 -460
rect 1760 -520 1780 -480
rect 1780 -520 1820 -480
rect 1820 -520 1840 -480
rect 5560 -40 5640 40
rect 1760 -540 1840 -520
rect 1220 -1040 1300 -960
rect 2220 -1100 2420 -900
rect 2960 -1100 3160 -900
rect 4360 -880 4440 -860
rect 4360 -920 4380 -880
rect 4380 -920 4420 -880
rect 4420 -920 4440 -880
rect 4360 -940 4440 -920
rect 2280 -1340 2360 -1260
rect 5920 -920 6120 -900
rect 5920 -1080 5980 -920
rect 5980 -1080 6060 -920
rect 6060 -1080 6120 -920
rect 5920 -1100 6120 -1080
rect 1580 -1760 1660 -1680
rect 3480 -2020 3560 -1940
rect 1820 -2330 1900 -2320
rect 1900 -2330 1940 -2320
rect 1940 -2330 2020 -2320
rect 1820 -2520 2020 -2330
rect 1120 -2820 1200 -2740
rect 4400 -2940 4600 -2740
rect 3000 -3080 3080 -3060
rect 3000 -3120 3020 -3080
rect 3020 -3120 3060 -3080
rect 3060 -3120 3080 -3080
rect 3000 -3140 3080 -3120
rect 6620 -1760 6720 -1660
rect 6360 -1900 6440 -1820
rect 4980 -2920 5140 -2760
rect 360 -3420 560 -3220
rect 780 -3950 860 -3870
rect 3000 -4100 3120 -3960
rect 3000 -4140 3020 -4100
rect 3020 -4140 3060 -4100
rect 3060 -4140 3120 -4100
rect 3000 -4180 3120 -4140
<< metal2 >>
rect 3240 4160 3440 4166
rect 1160 3840 2280 3920
rect 2360 3840 2366 3920
rect 1160 2040 1240 3840
rect 3240 3640 3440 3960
rect 3240 3560 3300 3640
rect 3380 3560 3440 3640
rect 1580 3440 1780 3446
rect 1154 1960 1160 2040
rect 1240 1960 1540 2040
rect 660 780 780 800
rect 660 700 680 780
rect 760 700 1260 780
rect 1340 700 1346 780
rect 660 680 780 700
rect 360 100 980 300
rect 1180 100 1186 300
rect 360 -2320 560 100
rect 660 -960 780 -940
rect 660 -1040 680 -960
rect 760 -1040 1220 -960
rect 1300 -1040 1306 -960
rect 660 -1060 780 -1040
rect 1460 -1680 1540 1960
rect 1580 940 1780 3240
rect 2654 1080 2660 1160
rect 2740 1080 2746 1160
rect 1580 860 1620 940
rect 1740 860 1780 940
rect 1580 -380 1780 860
rect 1580 -460 2420 -380
rect 1580 -540 1760 -460
rect 1840 -540 2420 -460
rect 1580 -580 2420 -540
rect 2220 -900 2420 -580
rect 2220 -1260 2420 -1100
rect 2220 -1340 2280 -1260
rect 2360 -1340 2420 -1260
rect 2220 -1400 2420 -1340
rect 1580 -1680 1660 -1674
rect 1460 -1760 1580 -1680
rect 1580 -1766 1660 -1760
rect 360 -2520 1820 -2320
rect 2020 -2520 2026 -2320
rect 360 -3220 560 -2520
rect 2660 -2740 2740 1080
rect 3240 1040 3440 3560
rect 4960 2440 5080 2460
rect 3574 2360 3580 2440
rect 3660 2360 4980 2440
rect 5060 2360 5080 2440
rect 4960 2340 5080 2360
rect 3240 980 4900 1040
rect 3240 900 3300 980
rect 3380 900 4900 980
rect 3240 840 4900 900
rect 2800 300 3000 306
rect 3240 300 3440 840
rect 4700 680 4900 840
rect 4700 600 4760 680
rect 4840 600 4900 680
rect 4760 594 4840 600
rect 3000 100 3440 300
rect 2800 94 3000 100
rect 5540 40 5660 60
rect 5540 -40 5560 40
rect 5640 -40 5660 40
rect 5540 -60 5660 -40
rect 4300 -860 4500 -800
rect 600 -2820 1120 -2740
rect 1200 -2820 2740 -2740
rect 2960 -900 3160 -894
rect 4300 -900 4360 -860
rect 3160 -940 4360 -900
rect 4440 -900 4500 -860
rect 4440 -940 5920 -900
rect 3160 -1100 5920 -940
rect 6120 -1100 6126 -900
rect 354 -3420 360 -3220
rect 560 -3420 566 -3220
rect 600 -3860 680 -2820
rect 2960 -3060 3160 -1100
rect 6600 -1660 6740 -1640
rect 6600 -1760 6620 -1660
rect 6720 -1760 6740 -1660
rect 6600 -1780 6740 -1760
rect 6360 -1820 6440 -1814
rect 6360 -1940 6440 -1900
rect 3474 -2020 3480 -1940
rect 3560 -2020 6440 -1940
rect 4960 -2330 5080 -2320
rect 6620 -2330 6720 -1780
rect 4960 -2340 6720 -2330
rect 4960 -2420 4980 -2340
rect 5060 -2420 6720 -2340
rect 4960 -2430 6720 -2420
rect 4960 -2440 5080 -2430
rect 4394 -2940 4400 -2740
rect 4600 -2760 5160 -2740
rect 4600 -2920 4980 -2760
rect 5140 -2920 5160 -2760
rect 4600 -2940 5160 -2920
rect 2960 -3140 3000 -3060
rect 3080 -3140 3160 -3060
rect 600 -3870 860 -3860
rect 600 -3950 780 -3870
rect 600 -3960 860 -3950
rect 2960 -3960 3160 -3140
rect 2960 -4180 3000 -3960
rect 3120 -4180 3160 -3960
rect 2960 -4220 3160 -4180
<< via2 >>
rect 680 700 760 780
rect 680 -1040 760 -960
rect 4980 2360 5060 2440
rect 5565 -35 5635 35
rect 4980 -2420 5060 -2340
rect 4980 -2920 5140 -2760
<< metal3 >>
rect 4960 2445 5080 2460
rect 4960 2355 4975 2445
rect 5065 2355 5080 2445
rect 4960 2340 5080 2355
rect 660 785 780 800
rect 660 695 675 785
rect 765 695 780 785
rect 660 680 780 695
rect 5540 39 5660 60
rect 5540 -39 5561 39
rect 5639 -39 5660 39
rect 5540 -60 5660 -39
rect 660 -955 780 -940
rect 660 -1045 675 -955
rect 765 -1045 780 -955
rect 660 -1060 780 -1045
rect 4960 -2335 5080 -2320
rect 4960 -2425 4975 -2335
rect 5065 -2425 5080 -2335
rect 4960 -2440 5080 -2425
rect 4960 -2760 5160 -2740
rect 4960 -2920 4980 -2760
rect 5140 -2920 5160 -2760
rect 4960 -2940 5160 -2920
<< via3 >>
rect 4975 2440 5065 2445
rect 4975 2360 4980 2440
rect 4980 2360 5060 2440
rect 5060 2360 5065 2440
rect 4975 2355 5065 2360
rect 675 780 765 785
rect 675 700 680 780
rect 680 700 760 780
rect 760 700 765 780
rect 675 695 765 700
rect 5561 35 5639 39
rect 5561 -35 5565 35
rect 5565 -35 5635 35
rect 5635 -35 5639 35
rect 5561 -39 5639 -35
rect 675 -960 765 -955
rect 675 -1040 680 -960
rect 680 -1040 760 -960
rect 760 -1040 765 -960
rect 675 -1045 765 -1040
rect 4975 -2340 5065 -2335
rect 4975 -2420 4980 -2340
rect 4980 -2420 5060 -2340
rect 5060 -2420 5065 -2340
rect 4975 -2425 5065 -2420
rect 4980 -2920 5140 -2760
<< metal4 >>
rect 4960 2445 5080 2460
rect 4960 2440 4975 2445
rect 4720 2360 4975 2440
rect 4960 2355 4975 2360
rect 5065 2355 5080 2445
rect 4960 2340 5080 2355
rect 660 785 780 800
rect 660 695 675 785
rect 765 780 780 785
rect 765 700 960 780
rect 765 695 780 700
rect 660 680 780 695
rect 5540 39 5660 60
rect 5540 -39 5561 39
rect 5639 -39 5660 39
rect 5540 -60 5660 -39
rect 5560 -320 5640 -60
rect 660 -955 780 -940
rect 660 -1045 675 -955
rect 765 -960 780 -955
rect 765 -1040 980 -960
rect 765 -1045 780 -1040
rect 660 -1060 780 -1045
rect 4960 -2335 5080 -2320
rect 4960 -2340 4975 -2335
rect 4700 -2420 4975 -2340
rect 4960 -2425 4975 -2420
rect 5065 -2425 5080 -2335
rect 4960 -2440 5080 -2425
rect 4960 -2760 5160 -2740
rect 4960 -2920 4980 -2760
rect 5140 -2780 5160 -2760
rect 5540 -2780 5660 -1500
rect 5140 -2900 5660 -2780
rect 5140 -2920 5160 -2900
rect 4960 -2940 5160 -2920
use sky130_fd_pr__cap_mim_m3_1_VCAG9S  XC1
timestamp 1769561617
transform 0 1 5600 -1 0 -900
box -686 -540 686 540
use sky130_fd_pr__cap_mim_m3_1_6QCY69  XCb
timestamp 1769561617
transform -1 0 2886 0 -1 2240
box -1986 -1840 1986 1840
use sky130_fd_pr__cap_mim_m3_1_6QCY69  XCbp
timestamp 1769561617
transform -1 0 2886 0 -1 -2160
box -1986 -1840 1986 1840
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM1
timestamp 1769561617
transform -1 0 4600 0 -1 358
box -278 -358 278 358
use sky130_fd_pr__pfet_g5v0d10v5_PGELCA  XM1p
timestamp 1769561617
transform -1 0 4600 0 -1 -582
box -308 -418 308 418
use sky130_fd_pr__nfet_g5v0d10v5_FJGQ2Y  XM2p
timestamp 1769561617
transform 1 0 6398 0 1 -1282
box -278 -758 278 758
use sky130_fd_pr__pfet_g5v0d10v5_KLP5N5  XM2
timestamp 1769561617
transform 0 1 3600 -1 0 2100
box -308 -1297 308 1297
use sky130_fd_pr__nfet_g5v0d10v5_FJGQ2Y  XM3
timestamp 1769561617
transform 0 1 3500 -1 0 600
box -278 -758 278 758
use sky130_fd_pr__pfet_g5v0d10v5_KLP5N5  XM3p
timestamp 1769561617
transform 0 1 3000 -1 0 -700
box -308 -1297 308 1297
use sky130_fd_pr__nfet_g5v0d10v5_J2FQJR  XM4
timestamp 1769561617
transform 0 1 3611 -1 0 3880
box -278 -1258 278 1258
use sky130_fd_pr__pfet_g5v0d10v5_E47KVH  XM4p
timestamp 1769561617
transform 0 -1 2900 1 0 -3910
box -308 -2297 308 2297
use sky130_fd_pr__nfet_g5v0d10v5_FJGQ2Y  XM5p
timestamp 1769561617
transform -1 0 6938 0 -1 -1282
box -278 -758 278 758
use sky130_fd_pr__pfet_g5v0d10v5_KLP5N5  XM5
timestamp 1769561617
transform 0 1 3600 -1 0 2700
box -308 -1297 308 1297
use sky130_fd_pr__nfet_g5v0d10v5_FJGQ2Y  XM6
timestamp 1769561617
transform 1 0 1200 0 1 1200
box -278 -758 278 758
use sky130_fd_pr__pfet_g5v0d10v5_KLP5N5  XM6p
timestamp 1769561617
transform -1 0 1160 0 -1 -1700
box -308 -1297 308 1297
use sky130_fd_pr__nfet_g5v0d10v5_J2FQJR  XM8
timestamp 1769561617
transform 0 1 3611 -1 0 3340
box -278 -1258 278 1258
use sky130_fd_pr__pfet_g5v0d10v5_E47KVH  XM8p
timestamp 1769561617
transform 0 -1 2900 1 0 -3310
box -308 -2297 308 2297
use sky130_fd_pr__nfet_g5v0d10v5_SMGAG4  XMa
timestamp 1769561617
transform 0 1 3050 -1 0 1140
box -278 -308 278 308
use sky130_fd_pr__pfet_g5v0d10v5_KLAZY6  XMap
timestamp 1769561617
transform 0 1 1920 -1 0 -1300
box -308 -397 308 397
use sky130_fd_pr__pfet_g5v0d10v5_7EJ6Y6  XMb
timestamp 1769561617
transform 0 -1 2100 1 0 1100
box -308 -547 308 547
use sky130_fd_pr__nfet_g5v0d10v5_6UEAUM  XMbp
timestamp 1769561617
transform 0 1 1920 -1 0 -2100
box -278 -383 278 383
use sky130_fd_pr__nfet_g5v0d10v5_FJGQ2Y  XMc
timestamp 1769561617
transform 0 1 4100 -1 0 1140
box -278 -758 278 758
use sky130_fd_pr__pfet_g5v0d10v5_KLP5N5  XMcp
timestamp 1769561617
transform 0 1 3600 -1 0 -1300
box -308 -1297 308 1297
<< labels >>
flabel metal1 1900 -1820 3560 -1780 0 FreeSans 1600 0 0 0 Yp
flabel space 4560 -2044 4600 -1620 0 FreeSans 1600 0 -1600 0 Xp
flabel metal2 760 -1040 1220 -960 0 FreeSans 1600 0 -4800 0 Qp
flabel metal1 2520 1260 2560 2100 0 FreeSans 1600 0 -1120 -480 Y
flabel metal1 4540 1740 4680 1780 0 FreeSans 1600 0 1600 -1600 X
flabel metal2 3660 2360 4980 2440 0 FreeSans 1600 0 6080 0 P
flabel metal2 1160 2040 1240 3920 0 FreeSans 1600 0 -1600 0 h
flabel metal2 1200 -2820 2740 -2740 0 FreeSans 1600 0 0 1600 t
flabel metal1 0 1900 200 2100 0 FreeSans 256 0 0 0 HLD
port 0 nsew
flabel metal1 0 -100 200 100 0 FreeSans 256 0 0 0 in
port 5 nsew
flabel metal1 0 -3900 200 -3700 0 FreeSans 256 0 0 0 VSS
port 3 nsew
flabel metal1 0 3700 200 3900 0 FreeSans 256 0 0 0 VDD
port 2 nsew
flabel via2 680 700 760 780 0 FreeSans 1600 0 -1600 0 Q
flabel metal1 0 -2900 200 -2700 0 FreeSans 256 0 0 0 TRK
port 1 nsew
flabel metal4 4980 -2420 5060 -2340 0 FreeSans 1600 0 0 0 Pp
flabel space 4640 -1700 6342 -1620 0 FreeSans 1600 0 0 1280 Xp
flabel metal1 4740 -3260 4820 -1620 0 FreeSans 1600 0 -1920 0 Xp
flabel metal1 7400 800 7600 1000 0 FreeSans 256 0 0 0 out
port 4 nsew
<< end >>
